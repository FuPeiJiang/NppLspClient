module scintilla

pub const invalid_position = -1
pub const sci_start = 2000
pub const sci_optional_start = 3000
pub const sci_lexer_start = 4000
pub const sci_addtext = 2001
pub const sci_addstyledtext = 2002
pub const sci_inserttext = 2003
pub const sci_changeinsertion = 2672
pub const sci_clearall = 2004
pub const sci_deleterange = 2645
pub const sci_cleardocumentstyle = 2005
pub const sci_getlength = 2006
pub const sci_getcharat = 2007
pub const sci_getcurrentpos = 2008
pub const sci_getanchor = 2009
pub const sci_getstyleat = 2010
pub const sci_redo = 2011
pub const sci_setundocollection = 2012
pub const sci_selectall = 2013
pub const sci_setsavepoint = 2014
pub const sci_getstyledtext = 2015
pub const sci_canredo = 2016
pub const sci_markerlinefromhandle = 2017
pub const sci_markerdeletehandle = 2018
pub const sci_getundocollection = 2019
pub const scws_invisible = 0
pub const scws_visiblealways = 1
pub const scws_visibleafterindent = 2
pub const scws_visibleonlyinindent = 3
pub const sci_getviewws = 2020
pub const sci_setviewws = 2021
pub const sctd_longarrow = 0
pub const sctd_strikeout = 1
pub const sci_gettabdrawmode = 2698
pub const sci_settabdrawmode = 2699
pub const sci_positionfrompoint = 2022
pub const sci_positionfrompointclose = 2023
pub const sci_gotoline = 2024
pub const sci_gotopos = 2025
pub const sci_setanchor = 2026
pub const sci_getcurline = 2027
pub const sci_getendstyled = 2028
pub const sc_eol_crlf = 0
pub const sc_eol_cr = 1
pub const sc_eol_lf = 2
pub const sci_converteols = 2029
pub const sci_geteolmode = 2030
pub const sci_seteolmode = 2031
pub const sci_startstyling = 2032
pub const sci_setstyling = 2033
pub const sci_getbuffereddraw = 2034
pub const sci_setbuffereddraw = 2035
pub const sci_settabwidth = 2036
pub const sci_gettabwidth = 2121
pub const sci_cleartabstops = 2675
pub const sci_addtabstop = 2676
pub const sci_getnexttabstop = 2677
pub const sc_cp_utf8 = 65001
pub const sci_setcodepage = 2037
pub const sc_ime_windowed = 0
pub const sc_ime_inline = 1
pub const sci_getimeinteraction = 2678
pub const sci_setimeinteraction = 2679
pub const marker_max = 31
pub const sc_mark_circle = 0
pub const sc_mark_roundrect = 1
pub const sc_mark_arrow = 2
pub const sc_mark_smallrect = 3
pub const sc_mark_shortarrow = 4
pub const sc_mark_empty = 5
pub const sc_mark_arrowdown = 6
pub const sc_mark_minus = 7
pub const sc_mark_plus = 8
pub const sc_mark_vline = 9
pub const sc_mark_lcorner = 10
pub const sc_mark_tcorner = 11
pub const sc_mark_boxplus = 12
pub const sc_mark_boxplusconnected = 13
pub const sc_mark_boxminus = 14
pub const sc_mark_boxminusconnected = 15
pub const sc_mark_lcornercurve = 16
pub const sc_mark_tcornercurve = 17
pub const sc_mark_circleplus = 18
pub const sc_mark_circleplusconnected = 19
pub const sc_mark_circleminus = 20
pub const sc_mark_circleminusconnected = 21
pub const sc_mark_background = 22
pub const sc_mark_dotdotdot = 23
pub const sc_mark_arrows = 24
pub const sc_mark_pixmap = 25
pub const sc_mark_fullrect = 26
pub const sc_mark_leftrect = 27
pub const sc_mark_available = 28
pub const sc_mark_underline = 29
pub const sc_mark_rgbaimage = 30
pub const sc_mark_bookmark = 31
pub const sc_mark_verticalbookmark = 32
pub const sc_mark_character = 10000
pub const sc_marknum_folderend = 25
pub const sc_marknum_folderopenmid = 26
pub const sc_marknum_foldermidtail = 27
pub const sc_marknum_foldertail = 28
pub const sc_marknum_foldersub = 29
pub const sc_marknum_folder = 30
pub const sc_marknum_folderopen = 31
pub const sc_mask_folders = u32(0xfe000000)
pub const sci_markerdefine = 2040
pub const sci_markersetfore = 2041
pub const sci_markersetback = 2042
pub const sci_markersetbackselected = 2292
pub const sci_markerenablehighlight = 2293
pub const sci_markeradd = 2043
pub const sci_markerdelete = 2044
pub const sci_markerdeleteall = 2045
pub const sci_markerget = 2046
pub const sci_markernext = 2047
pub const sci_markerprevious = 2048
pub const sci_markerdefinepixmap = 2049
pub const sci_markeraddset = 2466
pub const sci_markersetalpha = 2476
pub const sc_max_margin = 4
pub const sc_margin_symbol = 0
pub const sc_margin_number = 1
pub const sc_margin_back = 2
pub const sc_margin_fore = 3
pub const sc_margin_text = 4
pub const sc_margin_rtext = 5
pub const sc_margin_colour = 6
pub const sci_setmargintypen = 2240
pub const sci_getmargintypen = 2241
pub const sci_setmarginwidthn = 2242
pub const sci_getmarginwidthn = 2243
pub const sci_setmarginmaskn = 2244
pub const sci_getmarginmaskn = 2245
pub const sci_setmarginsensitiven = 2246
pub const sci_getmarginsensitiven = 2247
pub const sci_setmargincursorn = 2248
pub const sci_getmargincursorn = 2249
pub const sci_setmarginbackn = 2250
pub const sci_getmarginbackn = 2251
pub const sci_setmargins = 2252
pub const sci_getmargins = 2253
pub const style_default = 32
pub const style_linenumber = 33
pub const style_bracelight = 34
pub const style_bracebad = 35
pub const style_controlchar = 36
pub const style_indentguide = 37
pub const style_calltip = 38
pub const style_folddisplaytext = 39
pub const style_lastpredefined = 39
pub const style_max = 255
pub const sc_charset_ansi = 0
pub const sc_charset_default = 1
pub const sc_charset_baltic = 186
pub const sc_charset_chinesebig5 = 136
pub const sc_charset_easteurope = 238
pub const sc_charset_gb2312 = 134
pub const sc_charset_greek = 161
pub const sc_charset_hangul = 129
pub const sc_charset_mac = 77
pub const sc_charset_oem = 255
pub const sc_charset_russian = 204
pub const sc_charset_oem866 = 866
pub const sc_charset_cyrillic = 1251
pub const sc_charset_shiftjis = 128
pub const sc_charset_symbol = 2
pub const sc_charset_turkish = 162
pub const sc_charset_johab = 130
pub const sc_charset_hebrew = 177
pub const sc_charset_arabic = 178
pub const sc_charset_vietnamese = 163
pub const sc_charset_thai = 222
pub const sc_charset_8859_15 = 1000
pub const sci_styleclearall = 2050
pub const sci_stylesetfore = 2051
pub const sci_stylesetback = 2052
pub const sci_stylesetbold = 2053
pub const sci_stylesetitalic = 2054
pub const sci_stylesetsize = 2055
pub const sci_stylesetfont = 2056
pub const sci_styleseteolfilled = 2057
pub const sci_styleresetdefault = 2058
pub const sci_stylesetunderline = 2059
pub const sc_case_mixed = 0
pub const sc_case_upper = 1
pub const sc_case_lower = 2
pub const sc_case_camel = 3
pub const sci_stylegetfore = 2481
pub const sci_stylegetback = 2482
pub const sci_stylegetbold = 2483
pub const sci_stylegetitalic = 2484
pub const sci_stylegetsize = 2485
pub const sci_stylegetfont = 2486
pub const sci_stylegeteolfilled = 2487
pub const sci_stylegetunderline = 2488
pub const sci_stylegetcase = 2489
pub const sci_stylegetcharacterset = 2490
pub const sci_stylegetvisible = 2491
pub const sci_stylegetchangeable = 2492
pub const sci_stylegethotspot = 2493
pub const sci_stylesetcase = 2060
pub const sc_font_size_multiplier = 100
pub const sci_stylesetsizefractional = 2061
pub const sci_stylegetsizefractional = 2062
pub const sc_weight_normal = 400
pub const sc_weight_semibold = 600
pub const sc_weight_bold = 700
pub const sci_stylesetweight = 2063
pub const sci_stylegetweight = 2064
pub const sci_stylesetcharacterset = 2066
pub const sci_stylesethotspot = 2409
pub const sci_setselfore = 2067
pub const sci_setselback = 2068
pub const sci_getselalpha = 2477
pub const sci_setselalpha = 2478
pub const sci_getseleolfilled = 2479
pub const sci_setseleolfilled = 2480
pub const sci_setcaretfore = 2069
pub const sci_assigncmdkey = 2070
pub const sci_clearcmdkey = 2071
pub const sci_clearallcmdkeys = 2072
pub const sci_setstylingex = 2073
pub const sci_stylesetvisible = 2074
pub const sci_getcaretperiod = 2075
pub const sci_setcaretperiod = 2076
pub const sci_setwordchars = 2077
pub const sci_getwordchars = 2646
pub const sci_setcharactercategoryoptimization = 2720
pub const sci_getcharactercategoryoptimization = 2721
pub const sci_beginundoaction = 2078
pub const sci_endundoaction = 2079
pub const indic_plain = 0
pub const indic_squiggle = 1
pub const indic_tt = 2
pub const indic_diagonal = 3
pub const indic_strike = 4
pub const indic_hidden = 5
pub const indic_box = 6
pub const indic_roundbox = 7
pub const indic_straightbox = 8
pub const indic_dash = 9
pub const indic_dots = 10
pub const indic_squigglelow = 11
pub const indic_dotbox = 12
pub const indic_squigglepixmap = 13
pub const indic_compositionthick = 14
pub const indic_compositionthin = 15
pub const indic_fullbox = 16
pub const indic_textfore = 17
pub const indic_point = 18
pub const indic_pointcharacter = 19
pub const indic_gradient = 20
pub const indic_gradientcentre = 21
pub const indic_explorerlink = 22
pub const indic_container = 8
pub const indic_ime = 32
pub const indic_ime_max = 35
pub const indic_max = 35
pub const indicator_container = 8
pub const indicator_ime = 32
pub const indicator_ime_max = 35
pub const indicator_max = 35
pub const sci_indicsetstyle = 2080
pub const sci_indicgetstyle = 2081
pub const sci_indicsetfore = 2082
pub const sci_indicgetfore = 2083
pub const sci_indicsetunder = 2510
pub const sci_indicgetunder = 2511
pub const sci_indicsethoverstyle = 2680
pub const sci_indicgethoverstyle = 2681
pub const sci_indicsethoverfore = 2682
pub const sci_indicgethoverfore = 2683
pub const sc_indicvaluebit = 0x1000000
pub const sc_indicvaluemask = 0xffffff
pub const sc_indicflag_valuefore = 1
pub const sci_indicsetflags = 2684
pub const sci_indicgetflags = 2685
pub const sci_setwhitespacefore = 2084
pub const sci_setwhitespaceback = 2085
pub const sci_setwhitespacesize = 2086
pub const sci_getwhitespacesize = 2087
pub const sci_setlinestate = 2092
pub const sci_getlinestate = 2093
pub const sci_getmaxlinestate = 2094
pub const sci_getcaretlinevisible = 2095
pub const sci_setcaretlinevisible = 2096
pub const sci_getcaretlineback = 2097
pub const sci_setcaretlineback = 2098
pub const sci_getcaretlineframe = 2704
pub const sci_setcaretlineframe = 2705
pub const sci_stylesetchangeable = 2099
pub const sci_autocshow = 2100
pub const sci_autoccancel = 2101
pub const sci_autocactive = 2102
pub const sci_autocposstart = 2103
pub const sci_autoccomplete = 2104
pub const sci_autocstops = 2105
pub const sci_autocsetseparator = 2106
pub const sci_autocgetseparator = 2107
pub const sci_autocselect = 2108
pub const sci_autocsetcancelatstart = 2110
pub const sci_autocgetcancelatstart = 2111
pub const sci_autocsetfillups = 2112
pub const sci_autocsetchoosesingle = 2113
pub const sci_autocgetchoosesingle = 2114
pub const sci_autocsetignorecase = 2115
pub const sci_autocgetignorecase = 2116
pub const sci_userlistshow = 2117
pub const sci_autocsetautohide = 2118
pub const sci_autocgetautohide = 2119
pub const sci_autocsetdroprestofword = 2270
pub const sci_autocgetdroprestofword = 2271
pub const sci_registerimage = 2405
pub const sci_clearregisteredimages = 2408
pub const sci_autocgettypeseparator = 2285
pub const sci_autocsettypeseparator = 2286
pub const sci_autocsetmaxwidth = 2208
pub const sci_autocgetmaxwidth = 2209
pub const sci_autocsetmaxheight = 2210
pub const sci_autocgetmaxheight = 2211
pub const sci_setindent = 2122
pub const sci_getindent = 2123
pub const sci_setusetabs = 2124
pub const sci_getusetabs = 2125
pub const sci_setlineindentation = 2126
pub const sci_getlineindentation = 2127
pub const sci_getlineindentposition = 2128
pub const sci_getcolumn = 2129
pub const sci_countcharacters = 2633
pub const sci_countcodeunits = 2715
pub const sci_sethscrollbar = 2130
pub const sci_gethscrollbar = 2131
pub const sc_iv_none = 0
pub const sc_iv_real = 1
pub const sc_iv_lookforward = 2
pub const sc_iv_lookboth = 3
pub const sci_setindentationguides = 2132
pub const sci_getindentationguides = 2133
pub const sci_sethighlightguide = 2134
pub const sci_gethighlightguide = 2135
pub const sci_getlineendposition = 2136
pub const sci_getcodepage = 2137
pub const sci_getcaretfore = 2138
pub const sci_getreadonly = 2140
pub const sci_setcurrentpos = 2141
pub const sci_setselectionstart = 2142
pub const sci_getselectionstart = 2143
pub const sci_setselectionend = 2144
pub const sci_getselectionend = 2145
pub const sci_setemptyselection = 2556
pub const sci_setprintmagnification = 2146
pub const sci_getprintmagnification = 2147
pub const sc_print_normal = 0
pub const sc_print_invertlight = 1
pub const sc_print_blackonwhite = 2
pub const sc_print_colouronwhite = 3
pub const sc_print_colouronwhitedefaultbg = 4
pub const sc_print_screencolours = 5
pub const sci_setprintcolourmode = 2148
pub const sci_getprintcolourmode = 2149
pub const scfind_none = 0x0
pub const scfind_wholeword = 0x2
pub const scfind_matchcase = 0x4
pub const scfind_wordstart = 0x00100000
pub const scfind_regexp = 0x00200000
pub const scfind_posix = 0x00400000
pub const scfind_cxx11regex = 0x00800000
pub const sci_findtext = 2150
pub const sci_formatrange = 2151
pub const sci_getfirstvisibleline = 2152
pub const sci_getline = 2153
pub const sci_getlinecount = 2154
pub const sci_setmarginleft = 2155
pub const sci_getmarginleft = 2156
pub const sci_setmarginright = 2157
pub const sci_getmarginright = 2158
pub const sci_getmodify = 2159
pub const sci_setsel = 2160
pub const sci_getseltext = 2161
pub const sci_gettextrange = 2162
pub const sci_hideselection = 2163
pub const sci_pointxfromposition = 2164
pub const sci_pointyfromposition = 2165
pub const sci_linefromposition = 2166
pub const sci_positionfromline = 2167
pub const sci_linescroll = 2168
pub const sci_scrollcaret = 2169
pub const sci_scrollrange = 2569
pub const sci_replacesel = 2170
pub const sci_setreadonly = 2171
pub const sci_null = 2172
pub const sci_canpaste = 2173
pub const sci_canundo = 2174
pub const sci_emptyundobuffer = 2175
pub const sci_undo = 2176
pub const sci_cut = 2177
pub const sci_copy = 2178
pub const sci_paste = 2179
pub const sci_clear = 2180
pub const sci_settext = 2181
pub const sci_gettext = 2182
pub const sci_gettextlength = 2183
pub const sci_getdirectfunction = 2184
pub const sci_getdirectpointer = 2185
pub const sci_setovertype = 2186
pub const sci_getovertype = 2187
pub const sci_setcaretwidth = 2188
pub const sci_getcaretwidth = 2189
pub const sci_settargetstart = 2190
pub const sci_gettargetstart = 2191
pub const sci_settargetend = 2192
pub const sci_gettargetend = 2193
pub const sci_settargetrange = 2686
pub const sci_gettargettext = 2687
pub const sci_targetfromselection = 2287
pub const sci_targetwholedocument = 2690
pub const sci_replacetarget = 2194
pub const sci_replacetargetre = 2195
pub const sci_searchintarget = 2197
pub const sci_setsearchflags = 2198
pub const sci_getsearchflags = 2199
pub const sci_calltipshow = 2200
pub const sci_calltipcancel = 2201
pub const sci_calltipactive = 2202
pub const sci_calltipposstart = 2203
pub const sci_calltipsetposstart = 2214
pub const sci_calltipsethlt = 2204
pub const sci_calltipsetback = 2205
pub const sci_calltipsetfore = 2206
pub const sci_calltipsetforehlt = 2207
pub const sci_calltipusestyle = 2212
pub const sci_calltipsetposition = 2213
pub const sci_visiblefromdocline = 2220
pub const sci_doclinefromvisible = 2221
pub const sci_wrapcount = 2235
pub const sc_foldlevelbase = 0x400
pub const sc_foldlevelwhiteflag = 0x1000
pub const sc_foldlevelheaderflag = 0x2000
pub const sc_foldlevelnumbermask = 0x0fff
pub const sci_setfoldlevel = 2222
pub const sci_getfoldlevel = 2223
pub const sci_getlastchild = 2224
pub const sci_getfoldparent = 2225
pub const sci_showlines = 2226
pub const sci_hidelines = 2227
pub const sci_getlinevisible = 2228
pub const sci_getalllinesvisible = 2236
pub const sci_setfoldexpanded = 2229
pub const sci_getfoldexpanded = 2230
pub const sci_togglefold = 2231
pub const sci_togglefoldshowtext = 2700
pub const sc_folddisplaytext_hidden = 0
pub const sc_folddisplaytext_standard = 1
pub const sc_folddisplaytext_boxed = 2
pub const sci_folddisplaytextsetstyle = 2701
pub const sci_folddisplaytextgetstyle = 2707
pub const sci_setdefaultfolddisplaytext = 2722
pub const sci_getdefaultfolddisplaytext = 2723
pub const sc_foldaction_contract = 0
pub const sc_foldaction_expand = 1
pub const sc_foldaction_toggle = 2
pub const sci_foldline = 2237
pub const sci_foldchildren = 2238
pub const sci_expandchildren = 2239
pub const sci_foldall = 2662
pub const sci_ensurevisible = 2232
pub const sc_automaticfold_show = 0x0001
pub const sc_automaticfold_click = 0x0002
pub const sc_automaticfold_change = 0x0004
pub const sci_setautomaticfold = 2663
pub const sci_getautomaticfold = 2664
pub const sc_foldflag_linebefore_expanded = 0x0002
pub const sc_foldflag_linebefore_contracted = 0x0004
pub const sc_foldflag_lineafter_expanded = 0x0008
pub const sc_foldflag_lineafter_contracted = 0x0010
pub const sc_foldflag_levelnumbers = 0x0040
pub const sc_foldflag_linestate = 0x0080
pub const sci_setfoldflags = 2233
pub const sci_ensurevisibleenforcepolicy = 2234
pub const sci_settabindents = 2260
pub const sci_gettabindents = 2261
pub const sci_setbackspaceunindents = 2262
pub const sci_getbackspaceunindents = 2263
pub const sc_time_forever = 10000000
pub const sci_setmousedwelltime = 2264
pub const sci_getmousedwelltime = 2265
pub const sci_wordstartposition = 2266
pub const sci_wordendposition = 2267
pub const sci_israngeword = 2691
pub const sc_idlestyling_none = 0
pub const sc_idlestyling_tovisible = 1
pub const sc_idlestyling_aftervisible = 2
pub const sc_idlestyling_all = 3
pub const sci_setidlestyling = 2692
pub const sci_getidlestyling = 2693
pub const sc_wrap_none = 0
pub const sc_wrap_word = 1
pub const sc_wrap_char = 2
pub const sc_wrap_whitespace = 3
pub const sci_setwrapmode = 2268
pub const sci_getwrapmode = 2269
pub const sc_wrapvisualflag_none = 0x0000
pub const sc_wrapvisualflag_end = 0x0001
pub const sc_wrapvisualflag_start = 0x0002
pub const sc_wrapvisualflag_margin = 0x0004
pub const sci_setwrapvisualflags = 2460
pub const sci_getwrapvisualflags = 2461
pub const sc_wrapvisualflagloc_default = 0x0000
pub const sc_wrapvisualflagloc_end_by_text = 0x0001
pub const sc_wrapvisualflagloc_start_by_text = 0x0002
pub const sci_setwrapvisualflagslocation = 2462
pub const sci_getwrapvisualflagslocation = 2463
pub const sci_setwrapstartindent = 2464
pub const sci_getwrapstartindent = 2465
pub const sc_wrapindent_fixed = 0
pub const sc_wrapindent_same = 1
pub const sc_wrapindent_indent = 2
pub const sc_wrapindent_deepindent = 3
pub const sci_setwrapindentmode = 2472
pub const sci_getwrapindentmode = 2473
pub const sc_cache_none = 0
pub const sc_cache_caret = 1
pub const sc_cache_page = 2
pub const sc_cache_document = 3
pub const sci_setlayoutcache = 2272
pub const sci_getlayoutcache = 2273
pub const sci_setscrollwidth = 2274
pub const sci_getscrollwidth = 2275
pub const sci_setscrollwidthtracking = 2516
pub const sci_getscrollwidthtracking = 2517
pub const sci_textwidth = 2276
pub const sci_setendatlastline = 2277
pub const sci_getendatlastline = 2278
pub const sci_textheight = 2279
pub const sci_setvscrollbar = 2280
pub const sci_getvscrollbar = 2281
pub const sci_appendtext = 2282
pub const sc_phases_one = 0
pub const sc_phases_two = 1
pub const sc_phases_multiple = 2
pub const sci_getphasesdraw = 2673
pub const sci_setphasesdraw = 2674
pub const sc_eff_quality_mask = 0xf
pub const sc_eff_quality_default = 0
pub const sc_eff_quality_non_antialiased = 1
pub const sc_eff_quality_antialiased = 2
pub const sc_eff_quality_lcd_optimized = 3
pub const sci_setfontquality = 2611
pub const sci_getfontquality = 2612
pub const sci_setfirstvisibleline = 2613
pub const sc_multipaste_once = 0
pub const sc_multipaste_each = 1
pub const sci_setmultipaste = 2614
pub const sci_getmultipaste = 2615
pub const sci_gettag = 2616
pub const sci_linesjoin = 2288
pub const sci_linessplit = 2289
pub const sci_setfoldmargincolour = 2290
pub const sci_setfoldmarginhicolour = 2291
pub const sc_accessibility_disabled = 0
pub const sc_accessibility_enabled = 1
pub const sci_setaccessibility = 2702
pub const sci_getaccessibility = 2703
pub const sci_linedown = 2300
pub const sci_linedownextend = 2301
pub const sci_lineup = 2302
pub const sci_lineupextend = 2303
pub const sci_charleft = 2304
pub const sci_charleftextend = 2305
pub const sci_charright = 2306
pub const sci_charrightextend = 2307
pub const sci_wordleft = 2308
pub const sci_wordleftextend = 2309
pub const sci_wordright = 2310
pub const sci_wordrightextend = 2311
pub const sci_home = 2312
pub const sci_homeextend = 2313
pub const sci_lineend = 2314
pub const sci_lineendextend = 2315
pub const sci_documentstart = 2316
pub const sci_documentstartextend = 2317
pub const sci_documentend = 2318
pub const sci_documentendextend = 2319
pub const sci_pageup = 2320
pub const sci_pageupextend = 2321
pub const sci_pagedown = 2322
pub const sci_pagedownextend = 2323
pub const sci_edittoggleovertype = 2324
pub const sci_cancel = 2325
pub const sci_deleteback = 2326
pub const sci_tab = 2327
pub const sci_backtab = 2328
pub const sci_newline = 2329
pub const sci_formfeed = 2330
pub const sci_vchome = 2331
pub const sci_vchomeextend = 2332
pub const sci_zoomin = 2333
pub const sci_zoomout = 2334
pub const sci_delwordleft = 2335
pub const sci_delwordright = 2336
pub const sci_delwordrightend = 2518
pub const sci_linecut = 2337
pub const sci_linedelete = 2338
pub const sci_linetranspose = 2339
pub const sci_linereverse = 2354
pub const sci_lineduplicate = 2404
pub const sci_lowercase = 2340
pub const sci_uppercase = 2341
pub const sci_linescrolldown = 2342
pub const sci_linescrollup = 2343
pub const sci_deletebacknotline = 2344
pub const sci_homedisplay = 2345
pub const sci_homedisplayextend = 2346
pub const sci_lineenddisplay = 2347
pub const sci_lineenddisplayextend = 2348
pub const sci_homewrap = 2349
pub const sci_homewrapextend = 2450
pub const sci_lineendwrap = 2451
pub const sci_lineendwrapextend = 2452
pub const sci_vchomewrap = 2453
pub const sci_vchomewrapextend = 2454
pub const sci_linecopy = 2455
pub const sci_movecaretinsideview = 2401
pub const sci_linelength = 2350
pub const sci_bracehighlight = 2351
pub const sci_bracehighlightindicator = 2498
pub const sci_bracebadlight = 2352
pub const sci_bracebadlightindicator = 2499
pub const sci_bracematch = 2353
pub const sci_getvieweol = 2355
pub const sci_setvieweol = 2356
pub const sci_getdocpointer = 2357
pub const sci_setdocpointer = 2358
pub const sci_setmodeventmask = 2359
pub const edge_none = 0
pub const edge_line = 1
pub const edge_background = 2
pub const edge_multiline = 3
pub const sci_getedgecolumn = 2360
pub const sci_setedgecolumn = 2361
pub const sci_getedgemode = 2362
pub const sci_setedgemode = 2363
pub const sci_getedgecolour = 2364
pub const sci_setedgecolour = 2365
pub const sci_multiedgeaddline = 2694
pub const sci_multiedgeclearall = 2695
pub const sci_searchanchor = 2366
pub const sci_searchnext = 2367
pub const sci_searchprev = 2368
pub const sci_linesonscreen = 2370
pub const sc_popup_never = 0
pub const sc_popup_all = 1
pub const sc_popup_text = 2
pub const sci_usepopup = 2371
pub const sci_selectionisrectangle = 2372
pub const sci_setzoom = 2373
pub const sci_getzoom = 2374
pub const sc_documentoption_default = 0
pub const sc_documentoption_styles_none = 0x1
pub const sc_documentoption_text_large = 0x100
pub const sci_createdocument = 2375
pub const sci_addrefdocument = 2376
pub const sci_releasedocument = 2377
pub const sci_getdocumentoptions = 2379
pub const sci_getmodeventmask = 2378
pub const sci_setcommandevents = 2717
pub const sci_getcommandevents = 2718
pub const sci_setfocus = 2380
pub const sci_getfocus = 2381
pub const sc_status_ok = 0
pub const sc_status_failure = 1
pub const sc_status_badalloc = 2
pub const sc_status_warn_start = 1000
pub const sc_status_warn_regex = 1001
pub const sci_setstatus = 2382
pub const sci_getstatus = 2383
pub const sci_setmousedowncaptures = 2384
pub const sci_getmousedowncaptures = 2385
pub const sci_setmousewheelcaptures = 2696
pub const sci_getmousewheelcaptures = 2697
pub const sc_cursornormal = -1
pub const sc_cursorarrow = 2
pub const sc_cursorwait = 4
pub const sc_cursorreversearrow = 7
pub const sci_setcursor = 2386
pub const sci_getcursor = 2387
pub const sci_setcontrolcharsymbol = 2388
pub const sci_getcontrolcharsymbol = 2389
pub const sci_wordpartleft = 2390
pub const sci_wordpartleftextend = 2391
pub const sci_wordpartright = 2392
pub const sci_wordpartrightextend = 2393
pub const visible_slop = 0x01
pub const visible_strict = 0x04
pub const sci_setvisiblepolicy = 2394
pub const sci_dellineleft = 2395
pub const sci_dellineright = 2396
pub const sci_setxoffset = 2397
pub const sci_getxoffset = 2398
pub const sci_choosecaretx = 2399
pub const sci_grabfocus = 2400
pub const caret_slop = 0x01
pub const caret_strict = 0x04
pub const caret_jumps = 0x10
pub const caret_even = 0x08
pub const sci_setxcaretpolicy = 2402
pub const sci_setycaretpolicy = 2403
pub const sci_setprintwrapmode = 2406
pub const sci_getprintwrapmode = 2407
pub const sci_sethotspotactivefore = 2410
pub const sci_gethotspotactivefore = 2494
pub const sci_sethotspotactiveback = 2411
pub const sci_gethotspotactiveback = 2495
pub const sci_sethotspotactiveunderline = 2412
pub const sci_gethotspotactiveunderline = 2496
pub const sci_sethotspotsingleline = 2421
pub const sci_gethotspotsingleline = 2497
pub const sci_paradown = 2413
pub const sci_paradownextend = 2414
pub const sci_paraup = 2415
pub const sci_paraupextend = 2416
pub const sci_positionbefore = 2417
pub const sci_positionafter = 2418
pub const sci_positionrelative = 2670
pub const sci_positionrelativecodeunits = 2716
pub const sci_copyrange = 2419
pub const sci_copytext = 2420
pub const sc_sel_stream = 0
pub const sc_sel_rectangle = 1
pub const sc_sel_lines = 2
pub const sc_sel_thin = 3
pub const sci_setselectionmode = 2422
pub const sci_getselectionmode = 2423
pub const sci_getmoveextendsselection = 2706
pub const sci_getlineselstartposition = 2424
pub const sci_getlineselendposition = 2425
pub const sci_linedownrectextend = 2426
pub const sci_lineuprectextend = 2427
pub const sci_charleftrectextend = 2428
pub const sci_charrightrectextend = 2429
pub const sci_homerectextend = 2430
pub const sci_vchomerectextend = 2431
pub const sci_lineendrectextend = 2432
pub const sci_pageuprectextend = 2433
pub const sci_pagedownrectextend = 2434
pub const sci_stutteredpageup = 2435
pub const sci_stutteredpageupextend = 2436
pub const sci_stutteredpagedown = 2437
pub const sci_stutteredpagedownextend = 2438
pub const sci_wordleftend = 2439
pub const sci_wordleftendextend = 2440
pub const sci_wordrightend = 2441
pub const sci_wordrightendextend = 2442
pub const sci_setwhitespacechars = 2443
pub const sci_getwhitespacechars = 2647
pub const sci_setpunctuationchars = 2648
pub const sci_getpunctuationchars = 2649
pub const sci_setcharsdefault = 2444
pub const sci_autocgetcurrent = 2445
pub const sci_autocgetcurrenttext = 2610
pub const sc_caseinsensitivebehaviour_respectcase = 0
pub const sc_caseinsensitivebehaviour_ignorecase = 1
pub const sci_autocsetcaseinsensitivebehaviour = 2634
pub const sci_autocgetcaseinsensitivebehaviour = 2635
pub const sc_multiautoc_once = 0
pub const sc_multiautoc_each = 1
pub const sci_autocsetmulti = 2636
pub const sci_autocgetmulti = 2637
pub const sc_order_presorted = 0
pub const sc_order_performsort = 1
pub const sc_order_custom = 2
pub const sci_autocsetorder = 2660
pub const sci_autocgetorder = 2661
pub const sci_allocate = 2446
pub const sci_targetasutf8 = 2447
pub const sci_setlengthforencode = 2448
pub const sci_encodedfromutf8 = 2449
pub const sci_findcolumn = 2456
pub const sci_getcaretsticky = 2457
pub const sci_setcaretsticky = 2458
pub const sc_caretsticky_off = 0
pub const sc_caretsticky_on = 1
pub const sc_caretsticky_whitespace = 2
pub const sci_togglecaretsticky = 2459
pub const sci_setpasteconvertendings = 2467
pub const sci_getpasteconvertendings = 2468
pub const sci_selectionduplicate = 2469
pub const sc_alpha_transparent = 0
pub const sc_alpha_opaque = 255
pub const sc_alpha_noalpha = 256
pub const sci_setcaretlinebackalpha = 2470
pub const sci_getcaretlinebackalpha = 2471
pub const caretstyle_invisible = 0
pub const caretstyle_line = 1
pub const caretstyle_block = 2
pub const caretstyle_overstrike_bar = 0
pub const caretstyle_overstrike_block = 0x10
pub const caretstyle_ins_mask = 0xf
pub const caretstyle_block_after = 0x100
pub const sci_setcaretstyle = 2512
pub const sci_getcaretstyle = 2513
pub const sci_setindicatorcurrent = 2500
pub const sci_getindicatorcurrent = 2501
pub const sci_setindicatorvalue = 2502
pub const sci_getindicatorvalue = 2503
pub const sci_indicatorfillrange = 2504
pub const sci_indicatorclearrange = 2505
pub const sci_indicatorallonfor = 2506
pub const sci_indicatorvalueat = 2507
pub const sci_indicatorstart = 2508
pub const sci_indicatorend = 2509
pub const sci_setpositioncache = 2514
pub const sci_getpositioncache = 2515
pub const sci_copyallowline = 2519
pub const sci_getcharacterpointer = 2520
pub const sci_getrangepointer = 2643
pub const sci_getgapposition = 2644
pub const sci_indicsetalpha = 2523
pub const sci_indicgetalpha = 2524
pub const sci_indicsetoutlinealpha = 2558
pub const sci_indicgetoutlinealpha = 2559
pub const sci_setextraascent = 2525
pub const sci_getextraascent = 2526
pub const sci_setextradescent = 2527
pub const sci_getextradescent = 2528
pub const sci_markersymboldefined = 2529
pub const sci_marginsettext = 2530
pub const sci_margingettext = 2531
pub const sci_marginsetstyle = 2532
pub const sci_margingetstyle = 2533
pub const sci_marginsetstyles = 2534
pub const sci_margingetstyles = 2535
pub const sci_margintextclearall = 2536
pub const sci_marginsetstyleoffset = 2537
pub const sci_margingetstyleoffset = 2538
pub const sc_marginoption_none = 0
pub const sc_marginoption_sublineselect = 1
pub const sci_setmarginoptions = 2539
pub const sci_getmarginoptions = 2557
pub const sci_annotationsettext = 2540
pub const sci_annotationgettext = 2541
pub const sci_annotationsetstyle = 2542
pub const sci_annotationgetstyle = 2543
pub const sci_annotationsetstyles = 2544
pub const sci_annotationgetstyles = 2545
pub const sci_annotationgetlines = 2546
pub const sci_annotationclearall = 2547
pub const annotation_hidden = 0
pub const annotation_standard = 1
pub const annotation_boxed = 2
pub const annotation_indented = 3
pub const sci_annotationsetvisible = 2548
pub const sci_annotationgetvisible = 2549
pub const sci_annotationsetstyleoffset = 2550
pub const sci_annotationgetstyleoffset = 2551
pub const sci_releaseallextendedstyles = 2552
pub const sci_allocateextendedstyles = 2553
pub const undo_none = 0
pub const undo_may_coalesce = 1
pub const sci_addundoaction = 2560
pub const sci_charpositionfrompoint = 2561
pub const sci_charpositionfrompointclose = 2562
pub const sci_setmouseselectionrectangularswitch = 2668
pub const sci_getmouseselectionrectangularswitch = 2669
pub const sci_setmultipleselection = 2563
pub const sci_getmultipleselection = 2564
pub const sci_setadditionalselectiontyping = 2565
pub const sci_getadditionalselectiontyping = 2566
pub const sci_setadditionalcaretsblink = 2567
pub const sci_getadditionalcaretsblink = 2568
pub const sci_setadditionalcaretsvisible = 2608
pub const sci_getadditionalcaretsvisible = 2609
pub const sci_getselections = 2570
pub const sci_getselectionempty = 2650
pub const sci_clearselections = 2571
pub const sci_setselection = 2572
pub const sci_addselection = 2573
pub const sci_dropselectionn = 2671
pub const sci_setmainselection = 2574
pub const sci_getmainselection = 2575
pub const sci_setselectionncaret = 2576
pub const sci_getselectionncaret = 2577
pub const sci_setselectionnanchor = 2578
pub const sci_getselectionnanchor = 2579
pub const sci_setselectionncaretvirtualspace = 2580
pub const sci_getselectionncaretvirtualspace = 2581
pub const sci_setselectionnanchorvirtualspace = 2582
pub const sci_getselectionnanchorvirtualspace = 2583
pub const sci_setselectionnstart = 2584
pub const sci_getselectionnstart = 2585
pub const sci_setselectionnend = 2586
pub const sci_getselectionnend = 2587
pub const sci_setrectangularselectioncaret = 2588
pub const sci_getrectangularselectioncaret = 2589
pub const sci_setrectangularselectionanchor = 2590
pub const sci_getrectangularselectionanchor = 2591
pub const sci_setrectangularselectioncaretvirtualspace = 2592
pub const sci_getrectangularselectioncaretvirtualspace = 2593
pub const sci_setrectangularselectionanchorvirtualspace = 2594
pub const sci_getrectangularselectionanchorvirtualspace = 2595
pub const scvs_none = 0
pub const scvs_rectangularselection = 1
pub const scvs_useraccessible = 2
pub const scvs_nowraplinestart = 4
pub const sci_setvirtualspaceoptions = 2596
pub const sci_getvirtualspaceoptions = 2597
pub const sci_setrectangularselectionmodifier = 2598
pub const sci_getrectangularselectionmodifier = 2599
pub const sci_setadditionalselfore = 2600
pub const sci_setadditionalselback = 2601
pub const sci_setadditionalselalpha = 2602
pub const sci_getadditionalselalpha = 2603
pub const sci_setadditionalcaretfore = 2604
pub const sci_getadditionalcaretfore = 2605
pub const sci_rotateselection = 2606
pub const sci_swapmainanchorcaret = 2607
pub const sci_multipleselectaddnext = 2688
pub const sci_multipleselectaddeach = 2689
pub const sci_changelexerstate = 2617
pub const sci_contractedfoldnext = 2618
pub const sci_verticalcentrecaret = 2619
pub const sci_moveselectedlinesup = 2620
pub const sci_moveselectedlinesdown = 2621
pub const sci_setidentifier = 2622
pub const sci_getidentifier = 2623
pub const sci_rgbaimagesetwidth = 2624
pub const sci_rgbaimagesetheight = 2625
pub const sci_rgbaimagesetscale = 2651
pub const sci_markerdefinergbaimage = 2626
pub const sci_registerrgbaimage = 2627
pub const sci_scrolltostart = 2628
pub const sci_scrolltoend = 2629
pub const sc_technology_default = 0
pub const sc_technology_directwrite = 1
pub const sc_technology_directwriteretain = 2
pub const sc_technology_directwritedc = 3
pub const sci_settechnology = 2630
pub const sci_gettechnology = 2631
pub const sci_createloader = 2632
pub const sci_findindicatorshow = 2640
pub const sci_findindicatorflash = 2641
pub const sci_findindicatorhide = 2642
pub const sci_vchomedisplay = 2652
pub const sci_vchomedisplayextend = 2653
pub const sci_getcaretlinevisiblealways = 2654
pub const sci_setcaretlinevisiblealways = 2655
pub const sc_line_end_type_default = 0
pub const sc_line_end_type_unicode = 1
pub const sci_setlineendtypesallowed = 2656
pub const sci_getlineendtypesallowed = 2657
pub const sci_getlineendtypesactive = 2658
pub const sci_setrepresentation = 2665
pub const sci_getrepresentation = 2666
pub const sci_clearrepresentation = 2667

pub const sci_eolannotationsettext = 2740
pub const sci_eolannotationgettext = 2741
pub const sci_eolannotationsetstyle = 2742
pub const sci_eolannotationgetstyle = 2743
pub const sci_eolannotationclearall = 2744
pub const sci_eolannotationsetvisible = 2745
pub const sci_eolannotationgetvisible = 2746
pub const sci_eolannotationsetstyleoffset = 2747
pub const sci_eolannotationgetstyleoffset = 2748

pub const eolannotation_hidden = 0x0
pub const eolannotation_standard = 0x1
pub const eolannotation_boxed = 0x2
pub const eolannotation_stadium = 0x100
pub const eolannotation_flat_circle = 0x101
pub const eolannotation_angle_circle = 0x102
pub const eolannotation_circle_flat = 0x110
pub const eolannotation_flats = 0x111
pub const eolannotation_angle_flat = 0x112
pub const eolannotation_circle_angle = 0x120
pub const eolannotation_flat_angle = 0x121
pub const eolannotation_angles = 0x122

pub const sci_startrecord = 3001
pub const sci_stoprecord = 3002
pub const sci_setlexer = 4001
pub const sci_getlexer = 4002
pub const sci_colourise = 4003
pub const sci_setproperty = 4004

// keywordset_max 8
pub const keywordset_max = 30
pub const sci_setkeywords = 4005
pub const sci_setlexerlanguage = 4006
pub const sci_loadlexerlibrary = 4007
pub const sci_getproperty = 4008
pub const sci_getpropertyexpanded = 4009
pub const sci_getpropertyint = 4010
pub const sci_getlexerlanguage = 4012
pub const sci_privatelexercall = 4013
pub const sci_propertynames = 4014
pub const sc_type_boolean = 0
pub const sc_type_integer = 1
pub const sc_type_string = 2
pub const sci_propertytype = 4015
pub const sci_describeproperty = 4016
pub const sci_describekeywordsets = 4017
pub const sci_getlineendtypessupported = 4018
pub const sci_allocatesubstyles = 4020
pub const sci_getsubstylesstart = 4021
pub const sci_getsubstyleslength = 4022
pub const sci_getstylefromsubstyle = 4027
pub const sci_getprimarystylefromstyle = 4028
pub const sci_freesubstyles = 4023
pub const sci_setidentifiers = 4024
pub const sci_distancetosecondarystyles = 4025
pub const sci_getsubstylebases = 4026
pub const sci_getnamedstyles = 4029
pub const sci_nameofstyle = 4030
pub const sci_tagsofstyle = 4031
pub const sci_descriptionofstyle = 4032
pub const sc_mod_none = 0x0
pub const sc_mod_inserttext = 0x1
pub const sc_mod_deletetext = 0x2
pub const sc_mod_changestyle = 0x4
pub const sc_mod_changefold = 0x8
pub const sc_performed_user = 0x10
pub const sc_performed_undo = 0x20
pub const sc_performed_redo = 0x40
pub const sc_multistepundoredo = 0x80
pub const sc_laststepinundoredo = 0x100
pub const sc_mod_changemarker = 0x200
pub const sc_mod_beforeinsert = 0x400
pub const sc_mod_beforedelete = 0x800
pub const sc_multilineundoredo = 0x1000
pub const sc_startaction = 0x2000
pub const sc_mod_changeindicator = 0x4000
pub const sc_mod_changelinestate = 0x8000
pub const sc_mod_changemargin = 0x10000
pub const sc_mod_changeannotation = 0x20000
pub const sc_mod_container = 0x40000
pub const sc_mod_lexerstate = 0x80000
pub const sc_mod_insertcheck = 0x100000
pub const sc_mod_changetabstops = 0x200000
pub const sc_modeventmaskall = 0x3fffff
pub const sc_searchresult_linebuffermaxlength = 1024
pub const sc_update_content = 0x1
pub const sc_update_selection = 0x2
pub const sc_update_v_scroll = 0x4
pub const sc_update_h_scroll = 0x8
pub const scen_change = 768
pub const scen_setfocus = 512
pub const scen_killfocus = 256
pub const sck_down = 300
pub const sck_up = 301
pub const sck_left = 302
pub const sck_right = 303
pub const sck_home = 304
pub const sck_end = 305
pub const sck_prior = 306
pub const sck_next = 307
pub const sck_delete = 308
pub const sck_insert = 309
pub const sck_escape = 7
pub const sck_back = 8
pub const sck_tab = 9
pub const sck_return = 13
pub const sck_add = 310
pub const sck_subtract = 311
pub const sck_divide = 312
pub const sck_win = 313
pub const sck_rwin = 314
pub const sck_menu = 315
pub const scmod_norm = 0
pub const scmod_shift = 1
pub const scmod_ctrl = 2
pub const scmod_alt = 4
pub const scmod_super = 8
pub const scmod_meta = 16
pub const sc_ac_fillup = 1
pub const sc_ac_doubleclick = 2
pub const sc_ac_tab = 3
pub const sc_ac_newline = 4
pub const sc_ac_command = 5
pub const sc_charactersource_direct_input = 0
pub const sc_charactersource_tentative_input = 1
pub const sc_charactersource_ime_result = 2

pub const scn_styleneeded = 2000
pub const scn_charadded = 2001
pub const scn_savepointreached = 2002
pub const scn_savepointleft = 2003
pub const scn_modifyattemptro = 2004
pub const scn_key = 2005
pub const scn_doubleclick = 2006
pub const scn_updateui = 2007
pub const scn_modified = 2008
pub const scn_macrorecord = 2009
pub const scn_marginclick = 2010
pub const scn_needshown = 2011
pub const scn_painted = 2013
pub const scn_userlistselection = 2014
pub const scn_uridropped = 2015
pub const scn_dwellstart = 2016
pub const scn_dwellend = 2017
pub const scn_zoom = 2018
pub const scn_hotspotclick = 2019
pub const scn_hotspotdoubleclick = 2020
pub const scn_calltipclick = 2021
pub const scn_autocselection = 2022
pub const scn_indicatorclick = 2023
pub const scn_indicatorrelease = 2024
pub const scn_autoccancelled = 2025
pub const scn_autocchardeleted = 2026
pub const scn_hotspotreleaseclick = 2027
pub const scn_focusin = 2028
pub const scn_focusout = 2029
pub const scn_autoccompleted = 2030
pub const scn_marginrightclick = 2031
pub const scn_autocselectionchange = 2032

// provisional
pub const sc_bidirectional_disabled = 0
pub const sc_bidirectional_l2r = 1
pub const sc_bidirectional_r2l = 2
pub const sci_getbidirectional = 2708
pub const sci_setbidirectional = 2709
pub const sc_linecharacterindex_none = 0
pub const sc_linecharacterindex_utf32 = 1
pub const sc_linecharacterindex_utf16 = 2
pub const sci_getlinecharacterindex = 2710
pub const sci_allocatelinecharacterindex = 2711
pub const sci_releaselinecharacterindex = 2712
pub const sci_linefromindexposition = 2713
pub const sci_indexpositionfromline = 2714
